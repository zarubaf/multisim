../../axi/normal/src/cpu.sv