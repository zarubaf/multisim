../../normal/src/irq_loopback.sv