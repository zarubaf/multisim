../../normal/src/memory.sv