../../axi/normal/src/memory.sv