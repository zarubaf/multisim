../../normal/src/apb_pkg.sv