../../axi/normal/src/axi_pkg.sv